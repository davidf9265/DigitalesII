// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
// Created on Sat Oct 24 14:55:25 2009

// synthesis message_off 10175

`timescale 1ns/1ns

module N_N (
    reset,clock,S,CNT0,C,
    WA,WB,WR,DIRA0,DIRA1,DIRA2,DIRB0,DIRB1,DIRB2,DIRW0,DIRW1,DIRW2,EN_CNT,DIRRAM0,DIRRAM1,DIRRAM2,UD,LR,AS,RC,RIN,WIN,CLR,RRA,RRB,CM,DISTA,WC);

    input reset;
    input clock;
    input S;
    input CNT0;
    input C;
    tri0 reset;
    tri0 S;
    tri0 CNT0;
    tri0 C;
    output WA;
    output WB;
    output WR;
    output DIRA0;
    output DIRA1;
    output DIRA2;
    output DIRB0;
    output DIRB1;
    output DIRB2;
    output DIRW0;
    output DIRW1;
    output DIRW2;
    output EN_CNT;
    output DIRRAM0;
    output DIRRAM1;
    output DIRRAM2;
    output UD;
    output LR;
    output AS;
    output RC;
    output RIN;
    output WIN;
    output CLR;
    output RRA;
    output RRB;
    output CM;
    output DISTA;
    output WC;
    reg WA;
    reg WB;
    reg WR;
    reg DIRA0;
    reg DIRA1;
    reg DIRA2;
    reg DIRB0;
    reg DIRB1;
    reg DIRB2;
    reg DIRW0;
    reg DIRW1;
    reg DIRW2;
    reg EN_CNT;
    reg DIRRAM0;
    reg DIRRAM1;
    reg DIRRAM2;
    reg UD;
    reg LR;
    reg AS;
    reg RC;
    reg RIN;
    reg WIN;
    reg CLR;
    reg RRA;
    reg RRB;
    reg CM;
    reg DISTA;
    reg WC;
    reg [18:0] fstate;
    reg [18:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4,state6=5,state7=6,state8=7,state10=8,state11=9,state12=10,state13=11,state14=12,state15=13,state16=14,state17=15,state18=16,state9=17,state19=18;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or S or CNT0 or C)
    begin
        if (reset) begin
            reg_fstate <= state1;
            WA <= 1'b0;
            WB <= 1'b0;
            WR <= 1'b0;
            DIRA0 <= 1'b0;
            DIRA1 <= 1'b0;
            DIRA2 <= 1'b0;
            DIRB0 <= 1'b0;
            DIRB1 <= 1'b0;
            DIRB2 <= 1'b0;
            DIRW0 <= 1'b0;
            DIRW1 <= 1'b0;
            DIRW2 <= 1'b0;
            EN_CNT <= 1'b0;
            DIRRAM0 <= 1'b0;
            DIRRAM1 <= 1'b0;
            DIRRAM2 <= 1'b0;
            UD <= 1'b0;
            LR <= 1'b0;
            AS <= 1'b0;
            RC <= 1'b0;
            RIN <= 1'b0;
            WIN <= 1'b0;
            CLR <= 1'b0;
            RRA <= 1'b0;
            RRB <= 1'b0;
            CM <= 1'b0;
            DISTA <= 1'b0;
            WC <= 1'b0;
        end
        else begin
            WA <= 1'b0;
            WB <= 1'b0;
            WR <= 1'b0;
            DIRA0 <= 1'b0;
            DIRA1 <= 1'b0;
            DIRA2 <= 1'b0;
            DIRB0 <= 1'b0;
            DIRB1 <= 1'b0;
            DIRB2 <= 1'b0;
            DIRW0 <= 1'b0;
            DIRW1 <= 1'b0;
            DIRW2 <= 1'b0;
            EN_CNT <= 1'b0;
            DIRRAM0 <= 1'b0;
            DIRRAM1 <= 1'b0;
            DIRRAM2 <= 1'b0;
            UD <= 1'b0;
            LR <= 1'b0;
            AS <= 1'b0;
            RC <= 1'b0;
            RIN <= 1'b0;
            WIN <= 1'b0;
            CLR <= 1'b0;
            RRA <= 1'b0;
            RRB <= 1'b0;
            CM <= 1'b0;
            DISTA <= 1'b0;
            WC <= 1'b0;
            case (fstate)
                state1: begin
                    if (S)
                        reg_fstate <= state2;
                    else if (~(S))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    reg_fstate <= state19;

                    EN_CNT <= 1'b1;

                    DIRRAM0 <= 1'b1;

                    DIRRAM2 <= 1'b1;

                    CLR <= 1'b1;
                end
                state3: begin
                    if (CNT0)
                        reg_fstate <= state4;
                    else if (~(CNT0))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    EN_CNT <= 1'b1;

                    RIN <= 1'b1;

                    WIN <= 1'b1;

                    CM <= 1'b1;

                    WR <= 1'b1;
                end
                state4: begin
                    reg_fstate <= state5;

                    EN_CNT <= 1'b1;

                    UD <= 1'b1;
                end
                state5: begin
                    reg_fstate <= state6;

                    EN_CNT <= 1'b1;

                    DIRRAM1 <= 1'b0;

                    UD <= 1'b1;

                    DIRB0 <= 1'b1;

                    DIRB1 <= 1'b1;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA0 <= 1'b1;
                end
                state6: begin
                    reg_fstate <= state7;

                    DIRB0 <= 1'b1;

                    AS <= 1'b1;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    DISTA <= 1'b1;

                    WC <= 1'b1;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA1 <= 1'b1;
                end
                state7: begin
                    if (~(C))
                        reg_fstate <= state8;
                    else if (C)
                        reg_fstate <= state9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;
                end
                state8: begin
                    reg_fstate <= state5;

                    DIRW0 <= 1'b1;

                    RC <= 1'b1;

                    WR <= 1'b1;
                end
                state10: begin
                    if (C)
                        reg_fstate <= state11;
                    else if (~(C))
                        reg_fstate <= state13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state10;

                    EN_CNT <= 1'b0;

                    AS <= 1'b0;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    WC <= 1'b0;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA0 <= 1'b1;

                    DIRA2 <= 1'b1;
                end
                state11: begin
                    reg_fstate <= state12;

                    AS <= 1'b1;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    DISTA <= 1'b1;

                    WC <= 1'b1;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA0 <= 1'b1;
                end
                state12: begin
                    if (~(CNT0))
                        reg_fstate <= state17;
                    else if (CNT0)
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state12;

                    DIRW2 <= 1'b1;

                    DIRW0 <= 1'b1;

                    LR <= 1'b1;

                    AS <= 1'b1;

                    RC <= 1'b1;

                    DISTA <= 1'b1;

                    WC <= 1'b1;

                    WR <= 1'b1;
                end
                state13: begin
                    reg_fstate <= state14;

                    DIRW1 <= 1'b1;

                    AS <= 1'b1;

                    RC <= 1'b1;

                    RRA <= 1'b1;

                    DISTA <= 1'b1;

                    WC <= 1'b1;

                    WA <= 1'b1;

                    WR <= 1'b1;

                    DIRA2 <= 1'b1;
                end
                state14: begin
                    reg_fstate <= state15;

                    DIRW2 <= 1'b1;

                    DIRB2 <= 1'b0;

                    DIRW0 <= 1'b1;

                    RC <= 1'b1;

                    WR <= 1'b1;
                end
                state15: begin
                    reg_fstate <= state16;

                    DIRB0 <= 1'b1;

                    DIRB2 <= 1'b1;

                    RRB <= 1'b1;

                    WB <= 1'b1;
                end
                state16: begin
                    reg_fstate <= state12;

                    AS <= 1'b1;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    WC <= 1'b1;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA0 <= 1'b1;
                end
                state17: begin
                    reg_fstate <= state18;

                    DIRW0 <= 1'b1;

                    RC <= 1'b1;

                    WR <= 1'b1;
                end
                state18: begin
                    reg_fstate <= state9;

                    DIRB0 <= 1'b1;

                    RRA <= 1'b1;

                    RRB <= 1'b1;

                    WA <= 1'b1;

                    WB <= 1'b1;

                    DIRA1 <= 1'b1;
                end
                state9: begin
                    reg_fstate <= state10;

                    EN_CNT <= 1'b1;

                    AS <= 1'b0;

                    WC <= 1'b1;
                end
                state19: begin
                    reg_fstate <= state3;

                    EN_CNT <= 1'b1;

                    DIRRAM0 <= 1'b0;

                    DIRRAM2 <= 1'b1;

                    WIN <= 1'b1;
                end
                default: begin
                    WA <= 1'b0;
                    WB <= 1'b0;
                    WR <= 1'b0;
                    DIRA0 <= 1'b0;
                    DIRA1 <= 1'b0;
                    DIRA2 <= 1'b0;
                    DIRB0 <= 1'b0;
                    DIRB1 <= 1'b0;
                    DIRB2 <= 1'b0;
                    DIRW0 <= 1'b0;
                    DIRW1 <= 1'b0;
                    DIRW2 <= 1'b0;
                    EN_CNT <= 1'b0;
                    DIRRAM0 <= 1'b0;
                    DIRRAM1 <= 1'b0;
                    DIRRAM2 <= 1'b0;
                    UD <= 1'b0;
                    LR <= 1'b0;
                    AS <= 1'b0;
                    RC <= 1'b0;
                    RIN <= 1'b0;
                    WIN <= 1'b0;
                    CLR <= 1'b0;
                    RRA <= 1'b0;
                    RRB <= 1'b0;
                    CM <= 1'b0;
                    DISTA <= 1'b0;
                    WC <= 1'b0;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // N_N

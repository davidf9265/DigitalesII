-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 235 06/17/2009 Service Pack 2 SJ Web Edition
-- Created on Sat Oct 24 15:11:54 2009

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY N_N3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        S : IN STD_LOGIC := '0';
        CNT0 : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        WA : OUT STD_LOGIC;
        WB : OUT STD_LOGIC;
        WR : OUT STD_LOGIC;
        DIRA0 : OUT STD_LOGIC;
        DIRA1 : OUT STD_LOGIC;
        DIRA2 : OUT STD_LOGIC;
        DIRB0 : OUT STD_LOGIC;
        DIRB1 : OUT STD_LOGIC;
        DIRB2 : OUT STD_LOGIC;
        DIRW0 : OUT STD_LOGIC;
        DIRW1 : OUT STD_LOGIC;
        DIRW2 : OUT STD_LOGIC;
        EN_CNT : OUT STD_LOGIC;
        DIRRAM0 : OUT STD_LOGIC;
        DIRRAM1 : OUT STD_LOGIC;
        DIRRAM2 : OUT STD_LOGIC;
        UD : OUT STD_LOGIC;
        LR : OUT STD_LOGIC;
        AS : OUT STD_LOGIC;
        RC : OUT STD_LOGIC;
        RIN : OUT STD_LOGIC;
        WIN : OUT STD_LOGIC;
        CLR : OUT STD_LOGIC;
        RRA : OUT STD_LOGIC;
        RRB : OUT STD_LOGIC;
        CM : OUT STD_LOGIC;
        DISTA : OUT STD_LOGIC;
        WC : OUT STD_LOGIC
    );
END N_N3;

ARCHITECTURE BEHAVIOR OF N_N3 IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state8,state10,state11,state12,state13,state14,state15,state16,state17,state18,state19);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,S,CNT0,C)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            WA <= '0';
            WB <= '0';
            WR <= '0';
            DIRA0 <= '0';
            DIRA1 <= '0';
            DIRA2 <= '0';
            DIRB0 <= '0';
            DIRB1 <= '0';
            DIRB2 <= '0';
            DIRW0 <= '0';
            DIRW1 <= '0';
            DIRW2 <= '0';
            EN_CNT <= '0';
            DIRRAM0 <= '0';
            DIRRAM1 <= '0';
            DIRRAM2 <= '0';
            UD <= '0';
            LR <= '0';
            AS <= '0';
            RC <= '0';
            RIN <= '0';
            WIN <= '0';
            CLR <= '0';
            RRA <= '0';
            RRB <= '0';
            CM <= '0';
            DISTA <= '0';
            WC <= '0';
        ELSE
            WA <= '0';
            WB <= '0';
            WR <= '0';
            DIRA0 <= '0';
            DIRA1 <= '0';
            DIRA2 <= '0';
            DIRB0 <= '0';
            DIRB1 <= '0';
            DIRB2 <= '0';
            DIRW0 <= '0';
            DIRW1 <= '0';
            DIRW2 <= '0';
            EN_CNT <= '0';
            DIRRAM0 <= '0';
            DIRRAM1 <= '0';
            DIRRAM2 <= '0';
            UD <= '0';
            LR <= '0';
            AS <= '0';
            RC <= '0';
            RIN <= '0';
            WIN <= '0';
            CLR <= '0';
            RRA <= '0';
            RRB <= '0';
            CM <= '0';
            DISTA <= '0';
            WC <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF (NOT((S = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((S = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;
                WHEN state2 =>
                    reg_fstate <= state19;

                    EN_CNT <= '1';

                    DIRRAM2 <= '1';

                    DIRRAM0 <= '1';

                    CLR <= '1';
                WHEN state3 =>
                    IF ((CNT0 = '1')) THEN
                        reg_fstate <= state4;
                    ELSIF (NOT((CNT0 = '1'))) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    EN_CNT <= '1';

                    WIN <= '1';

                    RIN <= '1';

                    WR <= '1';

                    CM <= '1';
                WHEN state4 =>
                    reg_fstate <= state5;

                    UD <= '1';

                    EN_CNT <= '1';
                WHEN state5 =>
                    reg_fstate <= state6;

                    UD <= '1';

                    WA <= '1';

                    DIRB0 <= '1';

                    EN_CNT <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    DIRA0 <= '1';

                    DIRB1 <= '1';

                    WB <= '1';

                    DIRRAM1 <= '0';
                WHEN state6 =>
                    IF (NOT((C = '1'))) THEN
                        reg_fstate <= state8;
                    ELSIF ((C = '1')) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    WA <= '1';

                    DIRB0 <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    AS <= '1';

                    DIRA1 <= '1';

                    WB <= '1';

                    DISTA <= '1';

                    WC <= '1';
                WHEN state8 =>
                    reg_fstate <= state5;

                    RC <= '1';

                    DIRW0 <= '1';

                    WR <= '1';
                WHEN state10 =>
                    IF ((C = '1')) THEN
                        reg_fstate <= state11;
                    ELSIF (NOT((C = '1'))) THEN
                        reg_fstate <= state13;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    WA <= '1';

                    EN_CNT <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    DIRA0 <= '1';

                    WB <= '1';

                    DIRA2 <= '1';

                    WC <= '1';
                WHEN state11 =>
                    reg_fstate <= state12;

                    WA <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    DIRA0 <= '1';

                    AS <= '1';

                    WB <= '1';

                    DISTA <= '1';

                    WC <= '1';
                WHEN state12 =>
                    IF ((CNT0 = '1')) THEN
                        reg_fstate <= state1;
                    ELSIF (NOT((CNT0 = '1'))) THEN
                        reg_fstate <= state17;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state12;
                    END IF;

                    RC <= '1';

                    DIRW2 <= '1';

                    LR <= '1';

                    DIRW0 <= '1';

                    AS <= '1';

                    DISTA <= '1';

                    WR <= '1';

                    WC <= '1';
                WHEN state13 =>
                    reg_fstate <= state14;

                    WA <= '1';

                    RC <= '1';

                    RRA <= '1';

                    AS <= '1';

                    DIRA2 <= '1';

                    DISTA <= '1';

                    WR <= '1';

                    WC <= '1';

                    DIRW1 <= '1';
                WHEN state14 =>
                    reg_fstate <= state15;

                    RC <= '1';

                    DIRW2 <= '1';

                    DIRB2 <= '0';

                    DIRW0 <= '1';

                    WR <= '1';
                WHEN state15 =>
                    reg_fstate <= state16;

                    DIRB0 <= '1';

                    DIRB2 <= '1';

                    RRB <= '1';

                    WB <= '1';
                WHEN state16 =>
                    reg_fstate <= state12;

                    WA <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    DIRA0 <= '1';

                    AS <= '1';

                    WB <= '1';

                    WC <= '1';
                WHEN state17 =>
                    reg_fstate <= state18;

                    RC <= '1';

                    DIRW0 <= '1';

                    WR <= '1';
                WHEN state18 =>
                    reg_fstate <= state10;

                    WA <= '1';

                    DIRB0 <= '1';

                    RRB <= '1';

                    RRA <= '1';

                    DIRA1 <= '1';

                    WB <= '1';
                WHEN state19 =>
                    reg_fstate <= state3;

                    EN_CNT <= '1';

                    WIN <= '1';

                    DIRRAM2 <= '1';

                    DIRRAM0 <= '0';
                WHEN OTHERS => 
                    WA <= '0';
                    WB <= '0';
                    WR <= '0';
                    DIRA0 <= '0';
                    DIRA1 <= '0';
                    DIRA2 <= '0';
                    DIRB0 <= '0';
                    DIRB1 <= '0';
                    DIRB2 <= '0';
                    DIRW0 <= '0';
                    DIRW1 <= '0';
                    DIRW2 <= '0';
                    EN_CNT <= '0';
                    DIRRAM0 <= '0';
                    DIRRAM1 <= '0';
                    DIRRAM2 <= '0';
                    UD <= '0';
                    LR <= '0';
                    AS <= '0';
                    RC <= '0';
                    RIN <= '0';
                    WIN <= '0';
                    CLR <= '0';
                    RRA <= '0';
                    RRB <= '0';
                    CM <= '0';
                    DISTA <= '0';
                    WC <= '0';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
